`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12.11.2025 14:25:57
// Design Name: 
// Module Name: tb_half_adder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_half_adder(


    );
    reg a, b;
    wire sum, carry;
    half_adder uut(
    .a(a), .b(b), .sum(sum), .carry(carry)
    );
    initial begin
    a=0; b=0; #10;
    a=1; b=0; #10;
    a=0; b=1; #10;
    
endmodule
